module player_input (clk, reset, KEY, KEY_out);
	// This module is given a stabilized KEY input and outputs a pulse of the value.
	input logic 	clk, reset;
	input logic 	KEY;
	output logic 	KEY_out;
	enum { key_off, key_pulse, key_held } ps, ns;
	always_comb begin
			case (ps)
				key_off:		if (~KEY) 	ns = key_pulse;
								else			ns = key_off;
				key_pulse: 	if (~KEY) 	ns = key_held;
								else			ns = key_off;
				key_held: 	if (KEY)		ns = key_off;
								else 			ns = key_held;
			endcase
		end
	assign KEY_out = ps == key_pulse;
	always_ff @(posedge clk) begin
		if (reset)
			ps <= key_off;
		else
			ps <= ns;
	end
endmodule


module p_input_testbench();  
	 logic  clk, reset; 
	 logic  key;
	 logic  key_out;			
	  
	 p_input dut (clk, reset, key, key_out);   
		
	 // Set up a simulated clock.   
	 parameter CLOCK_PERIOD=100;  
	 initial begin  
	  clk <= 0;  
	  forever #(CLOCK_PERIOD/2) clk <= ~clk; // Forever toggle the clock 
	 end  
		
	 // Set up the inputs to the design.  Each line is a clock cycle.  
	 initial begin  
								 @(posedge clk);   
	  reset <= 1;         @(posedge clk); // Always reset FSMs at start  
	  reset <= 0; key <= 0; @(posedge clk);   
								 @(posedge clk);   
								 @(posedge clk);   
								 @(posedge clk);   
					  key <= 1; @(posedge clk);   
								 @(posedge clk);   
					  key <= 0; @(posedge clk);   
								 @(posedge clk);   
								 @(posedge clk);   
								 @(posedge clk);   
					  key <= 1; @(posedge clk);   
								 @(posedge clk);
					  reset <= 1;		 @(posedge clk); 
								 @(posedge clk); 
	  $stop; // End the simulation.  
	 end  
 endmodule